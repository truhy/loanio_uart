// soc_system.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                          //             clk.clk
		output wire        hps_0_h2f_reset_reset_n,          // hps_0_h2f_reset.reset_n
		output wire [66:0] hps_h2f_loan_io_in,               // hps_h2f_loan_io.in
		input  wire [66:0] hps_h2f_loan_io_out,              //                .out
		input  wire [66:0] hps_h2f_loan_io_oe,               //                .oe
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,  //          hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,    //                .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,    //                .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,    //                .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,    //                .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,    //                .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,    //                .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,     //                .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,  //                .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,  //                .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,  //                .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,    //                .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,    //                .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,    //                .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,      //                .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,       //                .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,       //                .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,      //                .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,       //                .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,       //                .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,       //                .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,       //                .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,       //                .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,       //                .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,       //                .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,       //                .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,       //                .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,       //                .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,      //                .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,      //                .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,      //                .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,      //                .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,     //                .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,    //                .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,    //                .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,     //                .hps_io_spim1_inst_SS0
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,      //                .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,      //                .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,      //                .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,      //                .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,   //                .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,   //                .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,   //                .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,   //                .hps_io_gpio_inst_GPIO61
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO49, //                .hps_io_gpio_inst_LOANIO49
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO50, //                .hps_io_gpio_inst_LOANIO50
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO53, //                .hps_io_gpio_inst_LOANIO53
		output wire [14:0] memory_mem_a,                     //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //                .mem_ba
		output wire        memory_mem_ck,                    //                .mem_ck
		output wire        memory_mem_ck_n,                  //                .mem_ck_n
		output wire        memory_mem_cke,                   //                .mem_cke
		output wire        memory_mem_cs_n,                  //                .mem_cs_n
		output wire        memory_mem_ras_n,                 //                .mem_ras_n
		output wire        memory_mem_cas_n,                 //                .mem_cas_n
		output wire        memory_mem_we_n,                  //                .mem_we_n
		output wire        memory_mem_reset_n,               //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                    //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                   //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                 //                .mem_dqs_n
		output wire        memory_mem_odt,                   //                .mem_odt
		output wire [3:0]  memory_mem_dm,                    //                .mem_dm
		input  wire        memory_oct_rzqin,                 //                .oct_rzqin
		input  wire        reset_reset_n                     //           reset.reset_n
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_loan_in               (hps_h2f_loan_io_in),               // h2f_loan_io.in
		.h2f_loan_out              (hps_h2f_loan_io_out),              //            .out
		.h2f_loan_oe               (hps_h2f_loan_io_oe),               //            .oe
		.mem_a                     (memory_mem_a),                     //      memory.mem_a
		.mem_ba                    (memory_mem_ba),                    //            .mem_ba
		.mem_ck                    (memory_mem_ck),                    //            .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                  //            .mem_ck_n
		.mem_cke                   (memory_mem_cke),                   //            .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                  //            .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                 //            .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                 //            .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                  //            .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),               //            .mem_reset_n
		.mem_dq                    (memory_mem_dq),                    //            .mem_dq
		.mem_dqs                   (memory_mem_dqs),                   //            .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                 //            .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                   //            .mem_odt
		.mem_dm                    (memory_mem_dm),                    //            .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                 //            .oct_rzqin
		.hps_io_emac1_inst_TX_CLK  (hps_io_hps_io_emac1_inst_TX_CLK),  //      hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0    (hps_io_hps_io_emac1_inst_TXD0),    //            .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1    (hps_io_hps_io_emac1_inst_TXD1),    //            .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2    (hps_io_hps_io_emac1_inst_TXD2),    //            .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3    (hps_io_hps_io_emac1_inst_TXD3),    //            .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0    (hps_io_hps_io_emac1_inst_RXD0),    //            .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO    (hps_io_hps_io_emac1_inst_MDIO),    //            .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC     (hps_io_hps_io_emac1_inst_MDC),     //            .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL  (hps_io_hps_io_emac1_inst_RX_CTL),  //            .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL  (hps_io_hps_io_emac1_inst_TX_CTL),  //            .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK  (hps_io_hps_io_emac1_inst_RX_CLK),  //            .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1    (hps_io_hps_io_emac1_inst_RXD1),    //            .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2    (hps_io_hps_io_emac1_inst_RXD2),    //            .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3    (hps_io_hps_io_emac1_inst_RXD3),    //            .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),      //            .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),       //            .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),       //            .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),      //            .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),       //            .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),       //            .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_io_hps_io_usb1_inst_D0),       //            .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_io_hps_io_usb1_inst_D1),       //            .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_io_hps_io_usb1_inst_D2),       //            .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_io_hps_io_usb1_inst_D3),       //            .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_io_hps_io_usb1_inst_D4),       //            .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_io_hps_io_usb1_inst_D5),       //            .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_io_hps_io_usb1_inst_D6),       //            .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_io_hps_io_usb1_inst_D7),       //            .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_io_hps_io_usb1_inst_CLK),      //            .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_io_hps_io_usb1_inst_STP),      //            .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_io_hps_io_usb1_inst_DIR),      //            .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_io_hps_io_usb1_inst_NXT),      //            .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK     (hps_io_hps_io_spim1_inst_CLK),     //            .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI    (hps_io_hps_io_spim1_inst_MOSI),    //            .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO    (hps_io_hps_io_spim1_inst_MISO),    //            .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0     (hps_io_hps_io_spim1_inst_SS0),     //            .hps_io_spim1_inst_SS0
		.hps_io_i2c0_inst_SDA      (hps_io_hps_io_i2c0_inst_SDA),      //            .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_io_hps_io_i2c0_inst_SCL),      //            .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA      (hps_io_hps_io_i2c1_inst_SDA),      //            .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL      (hps_io_hps_io_i2c1_inst_SCL),      //            .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09   (hps_io_hps_io_gpio_inst_GPIO09),   //            .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35   (hps_io_hps_io_gpio_inst_GPIO35),   //            .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO54   (hps_io_hps_io_gpio_inst_GPIO54),   //            .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61   (hps_io_hps_io_gpio_inst_GPIO61),   //            .hps_io_gpio_inst_GPIO61
		.hps_io_gpio_inst_LOANIO49 (hps_io_hps_io_gpio_inst_LOANIO49), //            .hps_io_gpio_inst_LOANIO49
		.hps_io_gpio_inst_LOANIO50 (hps_io_hps_io_gpio_inst_LOANIO50), //            .hps_io_gpio_inst_LOANIO50
		.hps_io_gpio_inst_LOANIO53 (hps_io_hps_io_gpio_inst_LOANIO53), //            .hps_io_gpio_inst_LOANIO53
		.h2f_rst_n                 (hps_0_h2f_reset_reset_n)           //   h2f_reset.reset_n
	);

endmodule
